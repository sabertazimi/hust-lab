/**
 * @module datapath
 * @brief data path, core of mips cpu
 */
module datapath
(
    
);
    
endmodule // datapath