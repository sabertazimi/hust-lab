`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// Company: Hust
// Engineer: sabertazimi
//
// Create Date: 2016/05/23 22:48:38
// Design Name: lab2
// Module Name: _4bit_to_7segment
// Project Name: verilog lab
// Target Devices: FPGA
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module _4bit_to_7segment(

    );
endmodule
