// `ifndef DEFINES_INCLUDED
// `define DEFINES_INCLUDED

`define ADD 0000
    
// `endif
