module _8leds(input [7:0] x_in, output [7:0] y_out);
	assign y_out = x_in;
endmodule