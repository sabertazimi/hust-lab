`timescale 1ns / 1ps

module _8leds_data(input [7:0] x_in, output [7:0] y_out);
	assign y_out = x_in;
endmodule
