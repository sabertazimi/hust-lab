`define ADD 0000
